library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_SIGNED.ALL;



entity registro_dividendo_B is
generic (n : natural := 8;
			m : natural := 4);
	port	(clk,	reset, load:	in std_logic;	
			 dividendo : in std_logic_vector(n - 1 downto 0);
			 salida : out std_logic_vector(n downto 0));

end registro_dividendo_B;

architecture Behavioral of registro_dividendo_B is

signal salidaAux : std_logic_vector(n downto 0);

begin

		
		

	PROCESS(clk,reset,load,dividendo,salidaAux)
		begin
			if reset = '1' then
				salidaAux <= (OTHERS => '0');
			elsif clk'event and clk = '1' then
				if load = '1' then
				salidaAux <= '0' & dividendo;
				end if;
			end if;
			salida <= salidaAux;
		end process;


end Behavioral;

